library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity game_controller_tb is
end game_controller_tb;


architecture testbench of game_controller_tb is



begin



end testbench;